ENTITY codificador IS
	PORT(t0, t1, t2, t3, t4, t5, t6, t7, t8, t9: IN BIT;
		  s: OUT BIT_VECTOR(3 DOWNTO 0));
END codificador;
-------------------------------------------------------------------------------------------------------------------------------------------------
ARCHITECTURE structural OF codificador IS
BEGIN
	