ENTITY demux1x4 IS
	PORT(