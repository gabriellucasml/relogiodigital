LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.std_logic_unsigned.ALL;

ENTITY dmux1xW IS
	GENERIC(W : NATURAL := 8;  --QUANTIDADE DE SAIDAS
			  V : NATURAL := 4); --TAMANHO DA PALAVRA BINARIA
	PORT(entrada : STD_LOGIC_VECTOR (V-1 DOWNTO 0);
	     